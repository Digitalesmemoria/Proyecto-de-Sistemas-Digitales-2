library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity controlador is
   port( 
			CLOCK: in std_logic;
			Reset: in std_logic;
			START: in std_logic;
			JUGAR: in std_logic;
			CONSULTAR: in std_logic;
			PRESIONO: in std_logic;
			REPETIDA: in std_logic;
			IGUAL_D1: in std_logic;
			IGUAL_D2: in std_logic;
			IGUAL_D3: in std_logic;
			IGUAL_D4: in std_logic;
			IGUAL_D5: in std_logic;
			IGUAL_D6: in std_logic;
			IGUAL_D7: in std_logic;
			IGUAL_D8: in std_logic;
			IGUAL_D9: in std_logic;
			IGUAL_D10: in std_logic;
			TIEMPO2: in std_logic;
			TIEMPO4: in std_logic;
			TIEMPO6: in std_logic;
			TIEMPO8: in std_logic;
			TIEMPO10: in std_logic;
			TIEMPO12: in std_logic;
			TIEMPO14: in std_logic;
			TIEMPO16: in std_logic;
			TIEMPO18: in std_logic;
			TIEMPO20: in std_logic;
			TIEMPO5: in std_logic;
			TIEMPO3: in std_logic;
			GUARDADO: in std_logic;
			EN_D1: OUT std_logic;
			EN_D2: OUT std_logic;
			EN_D3: OUT std_logic;
			EN_D4: OUT std_logic;
			EN_D5: OUT std_logic;
			EN_D6: OUT std_logic;
			EN_D7: OUT std_logic;
			EN_D8: OUT std_logic;
			EN_D9: OUT std_logic;
			EN_D10: OUT std_logic;
			EN_DATOIN: OUT std_logic;
			EN_FIGURA: OUT std_logic;
			CLC_FIGURA: OUT std_logic;
			EN_PUNTOS: OUT std_logic;
			CLC_PUNTOS: OUT std_logic;
			EN_MOSTRAR: OUT std_logic;
			CLC_MOSTRAR: OUT std_logic;
			EN_RELOJ: OUT std_logic;
			CLC_RELOJ: OUT std_logic;
			EN_RAM: OUT std_logic;
			W: OUT std_logic;
			MOSTRAR: OUT std_logic;
			GANO: OUT std_logic;
			PERDIO: OUT std_logic
			);
end controlador;



architecture COMPORTAMIENTO of controlador is
	TYPE estado IS (Ta,Tb,Tc,Td,Te,Tf,Tg,Th,Ti,Tj,Tk,Tl,Tm,Tn,Tp,Tq,Tr,Ts,Tt,Tu,Tv,Tw,Tx,Ty,Tz,Ta1,Tb1,Tc1,Td1,Te1,Tf1,Tg1,Th1,Ti1,Tj1,Tk1,Tl1,Tm1,Tn1,Tp1,Tq1,Tr1,Ts1,Tt1,Tu1,Tv1,Tw1,Tx1,Ty1,Tz1,Ta2,Tb2,Tc2,Td2,Te2,Tf2,Tg2,Th2,Ti2,Tj2,Tk2,Tl2,Tm2,Tn2,Tp2,Tq2,Tr2,Ts2,Tt2,Tu2,Tv2,Tw2,Tx2,Ty2,Tz2,Ta3,Tb3,Tc3,Td3,Te3,Tf3,Tg3,Th3,Ti3,Tj3,Tk3,Tl3,Tm3,Tn3,Tp3,Tq3,Tr3,Ts3,Tt3,Tu3,Tv3,Tw3,Tx3,Ty3,Tz3,Ta4,Tb4,Tc4,Td4,Te4,Tf4,Tg4,Th4,Ti4,Tj4,Tk4,Tl4,Tm4,Tn4,Tp4,Tq4,Tr4,Ts4,Tt4,Tu4,Tv4,Tw4,Tx4,Ty4,Tz4,Ta5,Tb5,Tc5,Td5,Te5,Tf5,Tg5,Th5,Ti5,Tj5,Tk5,Tl5,Tm5,Tn5,Tp5,Tq5,Tr5,Ts5,Tt5,Tu5,Tv5,Tw5,Tx5,Ty5,Tz5,Ta6,Tb6,Tc6,Td6,Te6,Tf6,Tg6,Th6,Ti6,Tj6,Tk6,Tl6,Tm6,Tn6,Tp6,Tq6,Tr6,Ts6,Tt6,Tu6,Tv6,Tw6,Tx6,Ty6,Tz6,Ta7,Tb7,Tc7,Td7,Te7,Tf7,Tg7,Th7,Ti7,Tj7,Tk7,Tl7,Tm7,Tn7,Tp7,Tq7,Tr7,Ts7,Tt7,Tu7,Tv7,Tw7,Tx7,Ty7,Tz7,Ta8,Tb8,Tc8,Td8,Te8,Tf8,Tg8,Th8,Ti8,Tj8,Tk8,Tl8,Tm8,Tn8,Tp8,Tq8,Tr8,Ts8,Tt8,Tu8,Tv8,Tw8,Tx8,Ty8,Tz8,Ta9,Tb9,Tc9,Td9,Te9,Tf9,Tg9,Th9,Ti9,Tj9,Tk9,Tl9,Tm9,Tn9,Tp9,Tq9,Tr9,Ts9,Tt9,Tu9);
	SIGNAL y : estado;
begin
 PROCESS (Reset,CLOCK)
 begin
	if Reset='0' then y<=Ta;
	elsif (CLOCK'event and Clock='1') then 
		case y is
			when Ta=> if (START='1') then y<=Tb; 
						 else y<=Ta;
						 end if;
			when Tb=> if (START='0') then y<=Tc; 
						 else y<=Tb;
						 end if;
			when Tc=> if (JUGAR='1') then y<=Td; 
						 else y<=Tc;
						 end if;
			when Td=> if (JUGAR='0') then y<=Te; 
						 else y<=Td;
						 end if;
			when Te=> y<=Tf;
			when Tf=> if (PRESIONO='1') then y<=Tg;
						 elsif (TIEMPO2='1') then y<=Tr9;	
						 else y<=Tf;
						 end if;
			when Tg=> if (PRESIONO='0') then y<=Th;
						 elsif (TIEMPO2='1') then y<=Tr9;	
						 else y<=Tg;
						 end if;
			when Th=> if (IGUAL_D1='1') then y<=Ti; 
						 else y<=Tr9;
						 end if;
			when Ti=> y<=Tj;
			when Tj=> if (REPETIDA='1') then y<=TJ; 
						 else y<=Tk;
						 end if;
			when Tk=> y<=Tl;
			when Tl=> if (PRESIONO='1') then y<=Tm;
						 elsif (TIEMPO4='1') then y<=Tr9;	
						 else y<=Tl;
						 end if;
			when Tm=> if (PRESIONO='0') then y<=Tn;
						 elsif (TIEMPO4='1') then y<=Tr9;	
						 else y<=Tm;
						 end if;
			when Tn=> if (IGUAL_D1='1') then y<=Tp; 
						 else y<=Tr9;
						 end if;
			when Tp=> y<=Tq;
			when Tq=> if (PRESIONO='1') then y<=Tr;
						 elsif (TIEMPO4='1') then y<=Tr9;	
						 else y<=Tq;
						 end if;
			when Tr=> if (PRESIONO='0') then y<=Ts;
						 elsif (TIEMPO4='1') then y<=Tr9;	
						 else y<=Tr;
						 end if;
			when Ts=> if (IGUAL_D2='1') then y<=Tt; 
						 else y<=Tr9;
						 end if;
			when Tt=> if (REPETIDA='1') then y<=Tt; 
						 else y<=Tu;
						 end if;
			when Tu=> y<=Tv;
			when Tv=> if (PRESIONO='1') then y<=Tw;
						 elsif (TIEMPO6='1') then y<=Tr9;	
						 else y<=Tv;
						 end if;
			when Tw=> if (PRESIONO='0') then y<=Tx;
						 elsif (TIEMPO6='1') then y<=Tr9;	
						 else y<=Tw;
						 end if;
			when Tx=> if (IGUAL_D1='1') then y<=Ty; 
						 else y<=Tr9;
						 end if;
			when Ty=> y<=Tz;
			when Tz=> if (PRESIONO='1') then y<=Ta1;
						 elsif (TIEMPO6='1') then y<=Tr9;	
						 else y<=Tz;
						 end if;
			when Ta1=> if (PRESIONO='0') then y<=Tb1;
						  elsif (TIEMPO6='1') then y<=Tr9;	
						  else y<=Ta1;
						  end if;
			when Tb1=> if (IGUAL_D2='1') then y<=Tc1; 
						 else y<=Tr9;
						 end if;
			when Tc1=> y<=Td1;
			when Td1=> if (PRESIONO='1') then y<=Te1;
						 elsif (TIEMPO6='1') then y<=Tr9;	
						 else y<=Td1;
						 end if;
			when Te1=> if (PRESIONO='0') then y<=Tf1;
						  elsif (TIEMPO6='1') then y<=Tr9;	
						  else y<=Te1;
						  end if;
			when Tf1=> if (IGUAL_D3='1') then y<=Tg1; 
						 else y<=Tr9;
						 end if;
			when Tg1=> if (REPETIDA='1') then y<=Tg1; 
						 else y<=Th1;
						 end if;
			when Th1=> y<=Ti1;
			when Ti1=> if (PRESIONO='1') then y<=Tj1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Ti1;
						 end if;
			when Tj1=> if (PRESIONO='0') then y<=Tk1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Tj1;
						 end if;
			when Tk1=> if (IGUAL_D1='1') then y<=Tl1; 
						 else y<=Tr9;
						 end if;
			when Tl1=> y<=Tm1;
			when Tm1=> if (PRESIONO='1') then y<=Tn1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Tm1;
						 end if;
			when Tn1=> if (PRESIONO='0') then y<=Tp1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Tn1;
						 end if;
			when Tp1=> if (IGUAL_D2='1') then y<=Tq1; 
						 else y<=Tr9;
						 end if;
			when Tq1=> y<=Tr1;
			when Tr1=> if (PRESIONO='1') then y<=Ts1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Tr1;
						 end if;
			when Ts1=> if (PRESIONO='0') then y<=Tt1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Ts1;
						 end if;
			when Tt1=>  if (IGUAL_D3='1') then y<=Tu1; 
						 else y<=Tr9;
						 end if;
			when Tu1=> y<=Tv1;
			when Tv1=> if (PRESIONO='1') then y<=Tw1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Tv1;
						 end if;
			when Tw1=> if (PRESIONO='0') then y<=Tx1;
						 elsif (TIEMPO8='1') then y<=Tr9;	
						 else y<=Tw1;
						 end if;
			when Tx1=>   if (IGUAL_D4='1') then y<=Ty1; 
						 else y<=Tr9;
						 end if;
			when Ty1=> if (REPETIDA='1') then y<=Ty1; 
						 else y<=Tz1;
						 end if;
			when Tz1=> y<=Ta2;
			when Ta2=> if (PRESIONO='1') then y<=Tb2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Ta2;
						 end if;
			when Tb2=> if (PRESIONO='0') then y<=Tc2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Tb2;
						 end if;
			when Tc2=> if (IGUAL_D1='1') then y<=Td2; 
						 else y<=Tr9;
						 end if;
			when Td2=> y<=Te2;
			when Te2=> if (PRESIONO='1') then y<=Tf2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Te2;
						 end if;
			when Tf2=> if (PRESIONO='0') then y<=Tg2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Tf2;
						 end if;
			when Tg2=>  if (IGUAL_D2='1') then y<=Th2; 
						 else y<=Tr9;
						 end if;
			when Th2=> y<=Ti2;
			when Ti2=> if (PRESIONO='1') then y<=Tj2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Ti2;
						 end if;
			when Tj2=> if (PRESIONO='0') then y<=Tk2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Tj2;
						 end if;
			when Tk2=> if (IGUAL_D3='1') then y<=Tl2; 
						 else y<=Tr9;
						 end if;
			when Tl2=> y<=Tm2;
			when Tm2=> if (PRESIONO='1') then y<=Tn2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Tm2;
						 end if;
			when Tn2=> if (PRESIONO='0') then y<=Tp2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Tn2;
						 end if;
			when Tp2=> if (IGUAL_D4='1') then y<=Tq2; 
						 else y<=Tr9;
						 end if;
			when Tq2=> y<=Tr2;
			when Tr2=> if (PRESIONO='1') then y<=Ts2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Tr2;
						 end if;
			when Ts2=> if (PRESIONO='0') then y<=Tt2;
						 elsif (TIEMPO10='1') then y<=Tr9;	
						 else y<=Ts2;
						 end if;
			when Tt2=>  if (IGUAL_D5='1') then y<=Tu2; 
						 else y<=Tr9;
						 end if;
			when Tu2=> if (REPETIDA='1') then y<=Tu2; 
						 else y<=Tv2;
						 end if;
			when Tv2=> y<=Tw2;
			when Tw2=>  if (PRESIONO='1') then y<=Tx2;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tw2;
						 end if;
			when Tx2=> if (PRESIONO='0') then y<=Ty2;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tx2;
						 end if;
			when Ty2=>  if (IGUAL_D1='1') then y<=Tz2; 
						 else y<=Tr9;
						 end if;
			when Tz2=> y<=Ta3;
			when Ta3=> if (PRESIONO='1') then y<=Tb3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Ta3;
						 end if;
			when Tb3=> if (PRESIONO='0') then y<=Tc3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tb3;
						 end if;
			when Tc3=> if (IGUAL_D2='1') then y<=Td3; 
						 else y<=Tr9;
						 end if;
			when Td3=> y<=Te3;
			when Te3=> if (PRESIONO='1') then y<=Tf3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Te3;
						 end if;
			when Tf3=> if (PRESIONO='0') then y<=Tg3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tf3;
						 end if;
			when Tg3=> if (IGUAL_D3='1') then y<=Th3; 
						 else y<=Tr9;
						 end if;
			when Th3=> y<=Ti3;
			when Ti3=> if (PRESIONO='1') then y<=Tj3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Ti3;
						 end if;
			when Tj3=> if (PRESIONO='0') then y<=Tk3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tj3;
						 end if;
			when Tk3=> if (IGUAL_D4='1') then y<=Tl3; 
						 else y<=Tr9;
						 end if;
			when Tl3=> y<=Tm3;
			when Tm3=> if (PRESIONO='1') then y<=Tn3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tm3;
						 end if;
			when Tn3=> if (PRESIONO='0') then y<=Tp3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tn3;
						 end if;
			when Tp3=> if (IGUAL_D5='1') then y<=Tq3; 
						 else y<=Tr9;
						 end if;
			when Tq3=> y<=Tr3; 
			when Tr3=>  if (PRESIONO='1') then y<=Ts3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Tr3;
						 end if;
			when Ts3=> if (PRESIONO='0') then y<=Tt3;
						 elsif (TIEMPO12='1') then y<=Tr9;	
						 else y<=Ts3;
						 end if;
			when Tt3=> if (IGUAL_D6='1') then y<=Tu3; 
						 else y<=Tr9;
						 end if;
			when Tu3=> if (REPETIDA='1') then y<=Tu3; 
						 else y<=Tv3;
						 end if;
			when Tv3=> y<=Tw3; 
			when Tw3=> if (PRESIONO='1') then y<=Tx3;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tw3;
						 end if;
			when Tx3=> if (PRESIONO='0') then y<=Ty3;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tx3;
						 end if;
			when Ty3=> if (IGUAL_D1='1') then y<=Tz3; 
						 else y<=Tr9;
						 end if; 
			when Tz3=> y<=Ta4; 
			when Ta4=> if (PRESIONO='1') then y<=Tb4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Ta4;
						 end if;
			when Tb4=> if (PRESIONO='0') then y<=Tc4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tb4;
						 end if;
			when Tc4=> if (IGUAL_D2='1') then y<=Td4; 
						 else y<=Tr9;
						 end if;
			when Td4=> y<=Te4; 
			when Te4=> if (PRESIONO='1') then y<=Tf4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Te4;
						 end if;
			when Tf4=> if (PRESIONO='0') then y<=Tg4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tf4;
						 end if;
			when Tg4=> if (IGUAL_D3='1') then y<=Th4; 
						 else y<=Tr9;
						 end if;
			when Th4=> y<=Ti4;
			when Ti4=> if (PRESIONO='1') then y<=Tj4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Ti4;
						 end if;
			when Tj4=> if (PRESIONO='0') then y<=Tk4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tj4;
						 end if;
			when Tk4=> if (IGUAL_D4='1') then y<=Tl4; 
						 else y<=Tr9;
						 end if;
			when Tl4=> y<=Tm4;
			when Tm4=> if (PRESIONO='1') then y<=Tn4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tm4;
						 end if;
			when Tn4=>  if (PRESIONO='0') then y<=Tp4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tn4;
						 end if;
			when Tp4=> if (IGUAL_D5='1') then y<=Tq4; 
						 else y<=Tr9;
						 end if;
			when Tq4=> y<=Tr4; 
			when Tr4=> if (PRESIONO='1') then y<=Ts4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tr4;
						 end if;
			when Ts4=> if (PRESIONO='0') then y<=Tt4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Ts4;
						 end if;
			when Tt4=> if (IGUAL_D6='1') then y<=Tu4; 
						 else y<=Tr9;
						 end if;
			when Tu4=> y<=Tv4; 
			when Tv4=> if (PRESIONO='1') then y<=Tw4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tv4;
						 end if;
			when Tw4=> if (PRESIONO='0') then y<=Tx4;
						 elsif (TIEMPO14='1') then y<=Tr9;	
						 else y<=Tw4;
						 end if;
			when Tx4=>  if (IGUAL_D7='1') then y<=Tu4; 
						 else y<=Tr9;
						 end if;
			when Ty4=> if (REPETIDA='1') then y<=Ty4; 
						 else y<=Tz4;
						 end if; 
			when Tz4=> y<=Ta5;
			when Ta5=> if (PRESIONO='1') then y<=Tb5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Ta5;
						 end if;
			when Tb5=> if (PRESIONO='0') then y<=Tc5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tb5;
						 end if;
			when Tc5=> if (IGUAL_D1='1') then y<=Td5; 
						 else y<=Tr9;
						 end if;
			when Td5=> y<=Te5;
			when Te5=> if (PRESIONO='1') then y<=Tf5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Te5;
						 end if;
			when Tf5=> if (PRESIONO='0') then y<=Tg5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tf5;
						 end if;
			when Tg5=> if (IGUAL_D2='1') then y<=Th5; 
						 else y<=Tr9;
						 end if;
			when Th5=> y<=Ti5;
			when Ti5=> if (PRESIONO='1') then y<=Tj5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Ti5;
						 end if;
			when Tj5=> if (PRESIONO='0') then y<=Tk5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tj5;
						 end if;
			when Tk5=> if (IGUAL_D3='1') then y<=Tl5; 
						 else y<=Tr9;
						 end if;
			when Tl5=> y<=Tm5;
			when Tm5=> if (PRESIONO='1') then y<=Tn5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tm5;
						 end if;
			when Tn5=> if (PRESIONO='0') then y<=Tp5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tn5;
						 end if;
			when Tp5=> if (IGUAL_D4='1') then y<=Tq5; 
						 else y<=Tr9;
						 end if;
			when Tq5=> y<=Tr5; 
			when Tr5=> if (PRESIONO='1') then y<=Ts5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tr5;
						 end if;
			when Ts5=> if (PRESIONO='0') then y<=Tt5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Ts5;
						 end if;
			when Tt5=> if (IGUAL_D5='1') then y<=Tu5; 
						 else y<=Tr9;
						 end if;
			when Tu5=> y<=Tv5;
			when Tv5=> if (PRESIONO='1') then y<=Tw5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tv5;
						 end if;
			when Tw5=> if (PRESIONO='0') then y<=Tx5;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tw5;
						 end if;
			when Tx5=> if (IGUAL_D6='1') then y<=Ty5; 
						 else y<=Tr9;
						 end if;
			when Ty5=> y<=Tz5; 
			when Tz5=> if (PRESIONO='1') then y<=Ta6;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Tz5;
						 end if;
			when Ta6=> if (PRESIONO='0') then y<=Tb6;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Ta6;
						 end if;
			when Tb6=>  if (IGUAL_D7='1') then y<=Tc6; 
						 else y<=Tr9;
						 end if;
			when Tc6=> y<=Td6;
			when Td6=> if (PRESIONO='1') then y<=Te6;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Td6;
						 end if;
			when Te6=> if (PRESIONO='0') then y<=Tf6;
						 elsif (TIEMPO16='1') then y<=Tr9;	
						 else y<=Te6;
						 end if;
			when Tf6=> if (IGUAL_D8='1') then y<=Tg6; 
						 else y<=Tr9;
						 end if;
			when Tg6=> if (REPETIDA='1') then y<=Tg6; 
						 else y<=Th6;
						 end if;
			when Th6=> y<=Ti6;
			when Ti6=> if (PRESIONO='1') then y<=Tj6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Ti6;
						 end if;
			when Tj6=> if (PRESIONO='0') then y<=Tk6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tj6;
						 end if;
			when Tk6=> if (IGUAL_D1='1') then y<=Tl6; 
						 else y<=Tr9;
						 end if;
			when Tl6=> y<=Tm6;
			when Tm6=>  if (PRESIONO='1') then y<=Tn6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tm6;
						 end if;
			when Tn6=> if (PRESIONO='0') then y<=Tp6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tn6;
						 end if;
			when Tp6=> if (IGUAL_D2='1') then y<=Tq6; 
						 else y<=Tr9;
						 end if;
			when Tq6=> y<=Tr6; 
			when Tr6=> if (PRESIONO='1') then y<=Ts6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tr6;
						 end if;
			when Ts6=> if (PRESIONO='0') then y<=Tt6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Ts6;
						 end if;
			when Tt6=> if (IGUAL_D3='1') then y<=Tu6; 
						 else y<=Tr9;
						 end if;
			when Tu6=> y<=Tv6;
			when Tv6=> if (PRESIONO='1') then y<=Tw6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tv6;
						 end if;
			when Tw6=>  if (PRESIONO='0') then y<=Tx6;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tw6;
						 end if;
			when Tx6=> if (IGUAL_D4='1') then y<=Ty6; 
						 else y<=Tr9;
						 end if;
			when Ty6=> y<=Tz6; 
			when Tz6=> if (PRESIONO='1') then y<=Ta7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tz6;
						 end if;
			when Ta7=> if (PRESIONO='0') then y<=Tb7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Ta7;
						 end if;
			when Tb7=> if (IGUAL_D5='1') then y<=Tc7; 
						 else y<=Tr9;
						 end if;
			when Tc7=> y<=Td7;
			when Td7=> if (PRESIONO='1') then y<=Te7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Td7;
						 end if;
			when Te7=> if (PRESIONO='0') then y<=Tf7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Te7;
						 end if;
			when Tf7=> if (IGUAL_D6='1') then y<=Tg7; 
						 else y<=Tr9;
						 end if;
			when Tg7=> y<=Th7;
			when Th7=> if (PRESIONO='1') then y<=Ti7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Th7;
						 end if;
			when Ti7=> if (PRESIONO='0') then y<=Tj7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Ti7;
						 end if;
			when Tj7=> if (IGUAL_D7='1') then y<=Tk7; 
						 else y<=Tr9;
						 end if;
			when Tk7=> y<=Tl7; 
			when Tl7=> if (PRESIONO='1') then y<=Tm7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tl7;
						 end if;
			when Tm7=> if (PRESIONO='0') then y<=Tn7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tm7;
						 end if;
			when Tn7=> if (IGUAL_D8='1') then y<=Tp7; 
						 else y<=Tr9;
						 end if;
			when Tp7=> y<=Tq7;
			when Tq7=> if (PRESIONO='1') then y<=Tr7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tq7;
						 end if;
			when Tr7=>  if (PRESIONO='0') then y<=Ts7;
						 elsif (TIEMPO18='1') then y<=Tr9;	
						 else y<=Tr7;
						 end if;
			when Ts7=> if (IGUAL_D9='1') then y<=Tt7; 
						 else y<=Tr9;
						 end if;
			when Tt7=> if (REPETIDA='1') then y<=Tt7; 
						 else y<=Tu7;
						 end if; 
			when Tu7=> y<=Tv7;
			when Tv7=> if (PRESIONO='1') then y<=Tw7;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tv7;
						 end if;
			when Tw7=> if (PRESIONO='0') then y<=Tx7;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tw7;
						 end if; 
			when Tx7=> if (IGUAL_D1='1') then y<=Ty7; 
						 else y<=Tr9;
						 end if;
			when Ty7=> y<=Tz7;
			when Tz7=>  if (PRESIONO='1') then y<=Ta8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tz7;
						 end if;
			when Ta8=> if (PRESIONO='0') then y<=Tb8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Ta8;
						 end if; 
			when Tb8=> if (IGUAL_D2='1') then y<=Tc8; 
						 else y<=Tr9;
						 end if;
			when Tc8=> y<=Td8;
			when Td8=> if (PRESIONO='1') then y<=Te8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Td8;
						 end if;
			when Te8=> if (PRESIONO='0') then y<=Tf8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Te8;
						 end if; 
			when Tf8=> if (IGUAL_D3='1') then y<=Tg8; 
						 else y<=Tr9;
						 end if;
			when Tg8=> y<=Th8;
			when Th8=> if (PRESIONO='1') then y<=Ti8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Th8;
						 end if;
			when Ti8=> if (PRESIONO='0') then y<=Tj8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Ti8;
						 end if; 
			when Tj8=> if (IGUAL_D4='1') then y<=Tk8; 
						 else y<=Tr9;
						 end if;
			when Tk8=> y<=Tl8;
			when Tl8=> if (PRESIONO='1') then y<=Tm8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tl8;
						 end if;
			when Tm8=> if (PRESIONO='0') then y<=Tn8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tm8;
						 end if; 
			when Tn8=> if (IGUAL_D5='1') then y<=Tp8; 
						 else y<=Tr9;
						 end if;
			when Tp8=> y<=Tq8;
			when Tq8=> if (PRESIONO='1') then y<=Tr8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tq8;
						 end if;
			when Tr8=> if (PRESIONO='0') then y<=Ts8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tr8;
						 end if; 
			when Ts8=> if (IGUAL_D6='1') then y<=Tt8; 
						 else y<=Tr9;
						 end if;
			when Tt8=> y<=Tu8;
			when Tu8=> if (PRESIONO='1') then y<=Tv8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tu8;
						 end if;
			when Tv8=> if (PRESIONO='0') then y<=Tw8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tv8;
						 end if;
			when Tw8=> if (IGUAL_D7='1') then y<=Tx8; 
						 else y<=Tr9;
						 end if;
			when Tx8=> y<=Ty8;
			when Ty8=> if (PRESIONO='1') then y<=Tz8;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Ty8;
						 end if; 
			when Tz8=>if (PRESIONO='0') then y<=Ta9;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tz8;
						 end if;
			when Ta9=> if (IGUAL_D8='1') then y<=Tb9; 
						 else y<=Tr9;
						 end if;
			when Tb9=> y<=Tc9; 
			when Tc9=>  if (PRESIONO='1') then y<=Td9;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tc9;
						 end if;
			when Td9=> if (PRESIONO='0') then y<=Te9;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Td9;
						 end if;
			when Te9=> if (IGUAL_D9='1') then y<=Tf9; 
						 else y<=Tr9;
						 end if; 
			when Tf9=> y<=Tg9; 
			when Tg9=> if (PRESIONO='1') then y<=Th9;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Tg9;
						 end if;
			when Th9=> if (PRESIONO='0') then y<=Ti9;
						 elsif (TIEMPO20='1') then y<=Tr9;	
						 else y<=Th9;
						 end if;
			when Ti9=> if (IGUAL_D10='1') then y<=Tj9; 
						 else y<=Tr9;
						 end if; 
			when Tj9=> y<=Tk9;
			when Tk9=> if (GUARDADO='1') then y<=Tl9; 
						 else y<=Tk9;
						 end if;
			when Tl9=> if (TIEMPO5='1') then y<=Tt9; 
						 else y<=Tl9;
						 end if;
			when Tt9=> y<=Tm9;
			when Tu9=> --------------------------------------- borrar
			when Tm9=> if (JUGAR='1') then y<=Td;
						 elsif (CONSULTAR='1') then y<=Tn9;	
						 else y<=Tm9;
						 end if; 
			when Tn9=> if (CONSULTAR='0') then y<=TP9; 
						 else y<=Tn9;
						 end if;
			when Tp9=> if (TIEMPO4='1') then y<=Tq9; 
						 else y<=Tp9;
						 end if;
			when Tq9=> y<=Tp9;
			when Tr9=> y<=Ts9; ---------Estado perdio
			when Ts9=> if (TIEMPO3='1') then y<=Tm9; 
						 else y<=Ts9;
						 end if;
		end case;
end if;
 END PROCESS;
PROCESS (y)
begin
		
			EN_D1<='0';
			EN_D2<='0';
			EN_D3<='0';
			EN_D4<='0';
			EN_D5<='0';
			EN_D6<='0';
			EN_D7<='0';
			EN_D8<='0';
			EN_D9<='0';
			EN_D10<='0';
			EN_DATOIN<='0';
			EN_FIGURA<='0';
			CLC_FIGURA<='0';
			EN_PUNTOS<='0';
			CLC_PUNTOS<='0';
			EN_MOSTRAR<='0';
			CLC_MOSTRAR<='0';
			EN_RELOJ<='0';
			CLC_RELOJ<='0';
			EN_RAM<='0';
			W<='0';
			MOSTRAR<='0';
			GANO<='0';
			PERDIO<='0';
		
		case y is
			when Ta=> CLC_FIGURA<='1'; CLC_PUNTOS<='1'; CLC_MOSTRAR<='1'; CLC_RELOJ<='1';
			when Tb=> 
			when Tc=> 
			when Td=> EN_FIGURA<='1';
			when Te=> 
			when Tf=> EN_RELOJ<='1';
			when Tg=> EN_RELOJ<='1';  EN_DATOIN<='1'; EN_D1<='1';
			when Th=> CLC_RELOJ<='1';
			when Ti=> EN_PUNTOS<='1';
			when Tj=> EN_FIGURA<='1';
			when Tk=> EN_D2<='1';
			when Tl=> EN_RELOJ<='1';
			when Tm=> EN_RELOJ<='1';  EN_DATOIN<='1';
			when Tn=> EN_RELOJ<='1';
			when Tp=> EN_PUNTOS<='1'; EN_RELOJ<='1';
			when Tq=> EN_RELOJ<='1';
			when Tr=> EN_RELOJ<='1';  EN_DATOIN<='1';
			when Ts=> CLC_RELOJ<='1'; 
					  if (IGUAL_D2='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Tt=> EN_FIGURA<='1';
			when Tu=> EN_D3<='1';	
			when Tv=> EN_RELOJ<='1'; 
			when Tw=> EN_RELOJ<='1';  EN_DATOIN<='1';
			when Tx=> EN_RELOJ<='1';
			when Ty=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tz=> EN_RELOJ<='1';
			when Ta1=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tb1=> EN_RELOJ<='1';
			when Tc1=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Td1=> EN_RELOJ<='1';
			when Te1=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tf1=> CLC_RELOJ<='1';
						if (IGUAL_D3='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Tg1=> EN_FIGURA<='1';
			when Th1=> EN_D4<='1';
			when Ti1=> EN_RELOJ<='1';
			when Tj1=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tk1=> EN_RELOJ<='1';
			when Tl1=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tm1=> EN_RELOJ<='1';
			when Tn1=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tp1=> EN_RELOJ<='1';
			when Tq1=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tr1=> EN_RELOJ<='1';
			when Ts1=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tt1=> EN_RELOJ<='1';
			when Tu1=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tv1=> EN_RELOJ<='1';
			when Tw1=> EN_DATOIN<='1'; EN_RELOJ<='1';					
			when Tx1=> CLC_RELOJ<='1';
					if (IGUAL_D4='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Ty1=> EN_FIGURA<='1';
			when Tz1=> EN_D5<='1';
			when Ta2=> EN_RELOJ<='1';
			when Tb2=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tc2=> EN_RELOJ<='1';
			when Td2=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Te2=> EN_RELOJ<='1';
			when Tf2=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tg2=> EN_RELOJ<='1';
			when Th2=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Ti2=> EN_RELOJ<='1';
			when Tj2=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tk2=> EN_RELOJ<='1';
			when Tl2=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tm2=> EN_RELOJ<='1';
			when Tn2=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tp2=> EN_RELOJ<='1';
			when Tq2=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tr2=> EN_RELOJ<='1';
			when Ts2=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tt2=> CLC_RELOJ<='1';
						if (IGUAL_D5='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Tu2=> EN_FIGURA<='1';
			when Tv2=> EN_D6<='1';
			when Tw2=> EN_RELOJ<='1';
			when Tx2=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Ty2=> EN_RELOJ<='1';
			when Tz2=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Ta3=> EN_RELOJ<='1';
			when Tb3=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tc3=> EN_RELOJ<='1';
			when Td3=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Te3=> EN_RELOJ<='1';
			when Tf3=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tg3=> EN_RELOJ<='1';
			when Th3=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Ti3=> EN_RELOJ<='1';
			when Tj3=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tk3=> EN_RELOJ<='1';
			when Tl3=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tm3=> EN_RELOJ<='1';
			when Tn3=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tp3=> EN_RELOJ<='1';
			when Tq3=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tr3=> EN_RELOJ<='1';
			when Ts3=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tt3=>  CLC_RELOJ<='1';
						if (IGUAL_D6='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Tu3=> EN_FIGURA<='1';
			when Tv3=> EN_D7<='1';
			when Tw3=> EN_RELOJ<='1';
			when Tx3=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Ty3=>  EN_RELOJ<='1';
			when Tz3=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Ta4=> EN_RELOJ<='1';
			when Tb4=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tc4=> EN_RELOJ<='1';
			when Td4=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Te4=> EN_RELOJ<='1';
			when Tf4=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tg4=> EN_RELOJ<='1';
			when Th4=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Ti4=> EN_RELOJ<='1';
			when Tj4=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tk4=> EN_RELOJ<='1';
			when Tl4=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tm4=> EN_RELOJ<='1';
			when Tn4=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tp4=> EN_RELOJ<='1';
			when Tq4=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tr4=> EN_RELOJ<='1';
			when Ts4=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tt4=> EN_RELOJ<='1';
			when Tu4=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tv4=> EN_RELOJ<='1';
			when Tw4=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tx4=> CLC_RELOJ<='1';
						if (IGUAL_D7='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Ty4=>  EN_FIGURA<='1';
			when Tz4=> EN_D8<='1';
			when Ta5=> EN_RELOJ<='1';
			when Tb5=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tc5=> EN_RELOJ<='1';
			when Td5=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Te5=> EN_RELOJ<='1';
			when Tf5=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tg5=> EN_RELOJ<='1';
			when Th5=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Ti5=> EN_RELOJ<='1';
			when Tj5=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tk5=> EN_RELOJ<='1';
			when Tl5=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tm5=> EN_RELOJ<='1';
			when Tn5=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tp5=> EN_RELOJ<='1';
			when Tq5=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tr5=> EN_RELOJ<='1';
			when Ts5=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tt5=> EN_RELOJ<='1';
			when Tu5=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tv5=> EN_RELOJ<='1';
			when Tw5=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tx5=> EN_RELOJ<='1';
			when Ty5=> EN_RELOJ<='1';
			when Tz5=> EN_RELOJ<='1';
			when Ta6=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tb6=> EN_RELOJ<='1';
			when Tc6=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Td6=> EN_RELOJ<='1';
			when Te6=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tf6=> CLC_RELOJ<='1';
						if (IGUAL_D8='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Tg6=> EN_FIGURA<='1';
			when Th6=> EN_D9<='1';
			when Ti6=> EN_RELOJ<='1';
			when Tj6=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tk6=> EN_RELOJ<='1';
			when Tl6=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tm6=> EN_RELOJ<='1';
			when Tn6=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tp6=> EN_RELOJ<='1';
			when Tq6=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tr6=> EN_RELOJ<='1';
			when Ts6=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tt6=> EN_RELOJ<='1';
			when Tu6=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tv6=> EN_RELOJ<='1';
			when Tw6=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tx6=> EN_RELOJ<='1';
			when Ty6=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tz6=>EN_RELOJ<='1';
			when Ta7=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tb7=> EN_RELOJ<='1';
			when Tc7=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Td7=> EN_RELOJ<='1';
			when Te7=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tf7=> EN_RELOJ<='1';
			when Tg7=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Th7=> EN_RELOJ<='1';
			when Ti7=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tj7=> EN_RELOJ<='1';
			when Tk7=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tl7=> EN_RELOJ<='1';
			when Tm7=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tn7=> EN_RELOJ<='1';
			when Tp7=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tq7=> EN_RELOJ<='1';
			when Tr7=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Ts7=>  CLC_RELOJ<='1';
						if (IGUAL_D9='1') then EN_PUNTOS<='1';
						 else EN_PUNTOS<='0';
						 end if;
			when Tt7=> EN_FIGURA<='1';
			when Tu7=> EN_D10<='1';
			when Tv7=> EN_RELOJ<='1';
			when Tw7=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tx7=> EN_RELOJ<='1';
			when Ty7=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tz7=> EN_RELOJ<='1';
			when Ta8=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tb8=> EN_RELOJ<='1';
			when Tc8=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Td8=> EN_RELOJ<='1';
			when Te8=> EN_DATOIN<='1';EN_RELOJ<='1';
			when Tf8=> EN_RELOJ<='1';
			when Tg8=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Th8=> EN_RELOJ<='1';
			when Ti8=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tj8=> EN_RELOJ<='1';
			when Tk8=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tl8=> EN_RELOJ<='1';
			when Tm8=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tn8=> EN_RELOJ<='1';
			when Tp8=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tq8=> EN_RELOJ<='1';
			when Tr8=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Ts8=> EN_RELOJ<='1';
			when Tt8=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tu8=> EN_RELOJ<='1';
			when Tv8=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Tw8=> EN_RELOJ<='1';
			when Tx8=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Ty8=>  EN_RELOJ<='1';
			when Tz8=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Ta9=> EN_RELOJ<='1';
			when Tb9=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tc9=> EN_RELOJ<='1';
			when Td9=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Te9=> EN_RELOJ<='1';
			when Tf9=> EN_RELOJ<='1'; EN_PUNTOS<='1';
			when Tg9=> EN_RELOJ<='1';
			when Th9=> EN_DATOIN<='1'; EN_RELOJ<='1';
			when Ti9=> CLC_RELOJ<='1';
			when Tj9=> EN_PUNTOS<='1';  
			when Tk9=> EN_RAM<='1'; W<='1';
			when Tl9=> EN_RELOJ<='1'; GANO<='1';
			when Tt9=> CLC_RELOJ<='1'; EN_MOSTRAR<='1';
			when Tm9=> CLC_FIGURA<='1'; CLC_PUNTOS<='1';  CLC_RELOJ<='1';
			when Tn9=> CLC_MOSTRAR<='1';
			when Tp9=> EN_RELOJ<='1'; MOSTRAR<='1';
			when Tq9=> EN_MOSTRAR<='1'; CLC_RELOJ<='1';
			when Tr9=> CLC_RELOJ<='1'; 
			when Ts9=> EN_RELOJ<='1'; PERDIO<='1';
			when Tu9=>
		end case;
 END PROCESS;
END COMPORTAMIENTO;


	
	
	
	
	
